//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/20/2024 05:26:12 PM
// Design Name: 
// Module Name: rh_file_pkg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


package rh_file_pkg;
    
    `timescale 1ns/1ps   
    `include "uvm_macros.svh"
    import uvm_pkg::*;  
    import top_pkg::*;
    import tlul_pkg::*; 
    import config_pkg::*;
    import iopmp_pkg::*; 

    localparam IOPMPNumChan           = 2;
    localparam IOPMPRegions           = 4;
       
    `include "uvm_transaction_rh.sv" 
    `include "uvm_sequence_rh.sv"       
                                                                                                                                
    `include "uvm_drv_rh.sv"             
    `include "uvm_mon_rh.sv"          
                                                                                                  
    `include "uvm_sco_rh.sv"                                
                            
    `include "uvm_agent_rh.sv"           
    `include "uvm_env_rh.sv"                          
                                                                                  
    `include "uvm_test_rh.sv"


endpackage