



`define HW_ZERO 1'b0
`define HW_ONE  1'b1
`define FULL_MODEL_M FULL_MODEL